module twiddle_w_value(
    input [2:0] index,
    output reg [23:0]  W_value
); //W 의 값의 LUT  

// 24비트중 상위 12비트는 실수 하위 12비트는 허수이다. 
// ex) 0.70711 이 실수인경우 부호있는 12비트 범위의 절대값의 최대값인 2048        x / 2048 = 0.70711 하고 계산하면 x = 0.70711 * 2048 = 1448 

always @ (*) begin
    case (index)
    3'b000 : begin
        W_value <= 24'h400000;          // (1 + j0) x/2048 = 1 ,  x = 2048, 정규화 - /2 1048 의 h - 400, 허수부분 - 0이므로 0
    end
    3'b001 : begin
        W_value <= 24'h3B2E78;          // 0.92388 + j(−0.38268), 실수부분 x = 0.92388 * 2048 / 2  946 의  h = 3b2, 허수부분 -0.38268 * 2048/2 = -0.392의 h = e78
    end
    3'b010 : begin
        W_value <= 24'h2D4D2C;          // 0.70711+j(−0.70711), 0.70711 * 1024 = 724 의 h = 2d4, -0.70711 * 1024 = -724 의 h = D2c
    end
    3'b011 : begin
        W_value <= 24'h188C4E;          // 0.38268+j(−0.92388) 0.38268 * 1024 =  392 의 h = 188, -0.92388 * 1024 = -946 의  h = c4e
    end
    3'b100 : begin
        W_value <= 24'h000C00;          // 0+j(−1)      -1*1024 = -1024 의 h = C00
    end
    3'b101 : begin
        W_value <= 24'hE78C4E;          // −0.38268+j(−0.92388) -0.38268 * 2048/2 = -0.392의 h = e78,  -0.92388 * 1024 = -946 의  h = c4e
    end
    3'b110 : begin
        W_value <= 24'hD2CD2C;          // −0.70711+j(−0.70711)  -0.70711 * 1024 = -724 의 h = D2c,   -0.70711 * 1024 = -724 의 h = D2c
    end
    3'b111 : begin
        W_value <= 24'hC4EE78;          // −0.92388+j(−0.38268)  -0.92388 * 1024 = -946 의  h = c4e, -0.38268 * 2048/2 = -0.392의 h = e78
    end
    endcase
end

endmodule